Declare ML Module "tacfork".

(** This module declare the fork tactic.

It can be used with the following syntax:

  tac >> f

where [tac] and [f] are two tactics. The first tactic [tac] is used to generate
a list of goals, and [f] is subsequently used to solve them, exactly as would do
[tac; first [solve [f] | idtac]]. There is a practical difference, though: the
tactic [f] is executed in a forked thread for each subgoal generated by [tac].

This will therefore badly fail on a system where [Unix.fork] is not disponible.

*)
